module digitub_scan(An,Digital,digout1,digout2,digout3,digout4);
input[7:0]An,Digital;
output[7:0]digout1,digout2,digout3,digout4;
assign digout2=
             (An[3:0]==4'h0)?7'b1000000:
             (An[3:0]==4'h1)?7'b1111001:
             (An[3:0]==4'h2)?7'b0100100:
             (An[3:0]==4'h3)?7'b0110000:
             (An[3:0]==4'h4)?7'b0011001:
             (An[3:0]==4'h5)?7'b0010010:
             (An[3:0]==4'h6)?7'b0000010:
             (An[3:0]==4'h7)?7'b1111000:
             (An[3:0]==4'h8)?7'b0000000:
             (An[3:0]==4'h9)?7'b0010000:
             (An[3:0]==4'hA)?7'b0001000:
             (An[3:0]==4'hB)?7'b0000011:
             (An[3:0]==4'hC)?7'b1000110:
             (An[3:0]==4'hD)?7'b0100001:
             (An[3:0]==4'hE)?7'b0000110:
             (An[3:0]==4'hF)?7'b0001110:7'b0;
assign digout3=
             (An[7:4]==4'h0)?7'b1000000:
             (An[7:4]==4'h1)?7'b1111001:
             (An[7:4]==4'h2)?7'b0100100:
             (An[7:4]==4'h3)?7'b0110000:
             (An[7:4]==4'h4)?7'b0011001:
             (An[7:4]==4'h5)?7'b0010010:
             (An[7:4]==4'h6)?7'b0000010:
             (An[7:4]==4'h7)?7'b1111000:
             (An[7:4]==4'h8)?7'b0000000:
             (An[7:4]==4'h9)?7'b0010000:
             (An[7:4]==4'hA)?7'b0001000:
             (An[7:4]==4'hB)?7'b0000011:
             (An[7:4]==4'hC)?7'b1000110:
             (An[7:4]==4'hD)?7'b0100001:
             (An[7:4]==4'hE)?7'b0000110:
             (An[7:4]==4'hF)?7'b0001110:7'b0;
assign digout4=
             (Digital[3:0]==4'h0)?7'b1000000:
             (Digital[3:0]==4'h1)?7'b1111001:
             (Digital[3:0]==4'h2)?7'b0100100:
             (Digital[3:0]==4'h3)?7'b0110000:
             (Digital[3:0]==4'h4)?7'b0011001:
             (Digital[3:0]==4'h5)?7'b0010010:
             (Digital[3:0]==4'h6)?7'b0000010:
             (Digital[3:0]==4'h7)?7'b1111000:
             (Digital[3:0]==4'h8)?7'b0000000:
             (Digital[3:0]==4'h9)?7'b0010000:
             (Digital[3:0]==4'hA)?7'b0001000:
             (Digital[3:0]==4'hB)?7'b0000011:
             (Digital[3:0]==4'hC)?7'b1000110:
             (Digital[3:0]==4'hD)?7'b0100001:
             (Digital[3:0]==4'hE)?7'b0000110:
             (Digital[3:0]==4'hF)?7'b0001110:7'b0;
assign digout1=
             (Digital[7:4]==4'h0)?7'b1000000:
             (Digital[7:4]==4'h1)?7'b1111001:
             (Digital[7:4]==4'h2)?7'b0100100:
             (Digital[7:4]==4'h3)?7'b0110000:
             (Digital[7:4]==4'h4)?7'b0011001:
             (Digital[7:4]==4'h5)?7'b0010010:
             (Digital[7:4]==4'h6)?7'b0000010:
             (Digital[7:4]==4'h7)?7'b1111000:
             (Digital[7:4]==4'h8)?7'b0000000:
             (Digital[7:4]==4'h9)?7'b0010000:
             (Digital[7:4]==4'hA)?7'b0001000:
             (Digital[7:4]==4'hB)?7'b0000011:
             (Digital[7:4]==4'hC)?7'b1000110:
             (Digital[7:4]==4'hD)?7'b0100001:
             (Digital[7:4]==4'hE)?7'b0000110:
             (Digital[7:4]==4'hF)?7'b0001110:7'b0;
				 endmodule
				 