module Pipeline_InsMem(reset,nop,PC_82,Ins);
input[6:0] PC_82;
input reset,nop;
output[31:0] Ins;
reg[31:0] Instruct;
assign Ins=nop? 32'b0:Instruct;//load-useð�շ�����nopΪ1��ֱ�ӽ�Ins��ֵΪ0

always@(*) 
 begin
	if(!reset) Instruct<=32'b0;
	else 
	 begin
		case(PC_82[6:0])
		 	 7'b0000000: Instruct<=32'b000010_00000000000000000001001101;     //j   reset
     7'b0000001: Instruct<=32'b000010_00000000000000000001010011;     //j   ILLOP
		 7'b0000010: Instruct<=32'b000000_11010_00000_00000_00000_001000; //jr  XADR
		 7'b0000011: Instruct<=32'b001001_00000_01000_0000000011000000; //addiu $t0, $zero, 192   0
		 7'b0000100: Instruct<=32'b101011_00000_01000_0000000000000000; //sw    $t0, 0($zero)
		 7'b0000101: Instruct<=32'b001001_00000_01000_0000000011111001; //addiu $t0, $zero, 249   1
		 7'b0000110: Instruct<=32'b101011_00000_01000_0000000000000100; //sw    $t0, 4($zero)
		 7'b0000111: Instruct<=32'b001001_00000_01000_0000000010100100; //addiu $t0, $zero, 164   2
		 7'b0001000: Instruct<=32'b101011_00000_01000_0000000000001000; //sw    $t0, 8($zero)
		 7'b0001001: Instruct<=32'b001001_00000_01000_0000000010110000; //addiu $t0, $zero, 176   3
		 7'b0001010: Instruct<=32'b101011_00000_01000_0000000000001100; //sw    $t0, 12($zero)
		 7'b0001011: Instruct<=32'b001001_00000_01000_0000000010011001; //addiu $t0, $zero, 153   4
		 7'b0001100: Instruct<=32'b101011_00000_01000_0000000000010000; //sw    $t0, 16($zero)
		 7'b0001101: Instruct<=32'b001001_00000_01000_0000000010010010; //addiu $t0, $zero, 146   5
		 7'b0001110: Instruct<=32'b101011_00000_01000_0000000000010100; //sw    $t0, 20($zero)
		 7'b0001111: Instruct<=32'b001001_00000_01000_0000000010000010; //addiu $t0, $zero, 130   6
		 7'b0010000: Instruct<=32'b101011_00000_01000_0000000000011000; //sw    $t0, 24($zero)
		 7'b0010001: Instruct<=32'b001001_00000_01000_0000000011111000; //addiu $t0, $zero, 248   7
		 7'b0010010: Instruct<=32'b101011_00000_01000_0000000000011100; //sw    $t0, 28($zero)
		 7'b0010011: Instruct<=32'b001001_00000_01000_0000000010000000; //addiu $t0, $zero, 128   8
		 7'b0010100: Instruct<=32'b101011_00000_01000_0000000000100000; //sw    $t0, 32($zero)
		 7'b0010101: Instruct<=32'b001001_00000_01000_0000000010010000; //addiu $t0, $zero, 144   9
		 7'b0010110: Instruct<=32'b101011_00000_01000_0000000000100100; //sw    $t0, 36($zero)
		 7'b0010111: Instruct<=32'b001001_00000_01000_0000000010001000; //addiu $t0, $zero, 136   a
		 7'b0011000: Instruct<=32'b101011_00000_01000_0000000000101000; //sw    $t0, 40($zero)
		 7'b0011001: Instruct<=32'b001001_00000_01000_0000000010000011; //addiu $t0, $zero, 131   b
		 7'b0011010: Instruct<=32'b101011_00000_01000_0000000000101100; //sw    $t0, 44($zero)
		 7'b0011011: Instruct<=32'b001001_00000_01000_0000000011000110; //addiu $t0, $zero, 198   c
		 7'b0011100: Instruct<=32'b101011_00000_01000_0000000000110000; //sw    $t0, 48$(zero)
		 7'b0011101: Instruct<=32'b001001_00000_01000_0000000010100001; //addiu $t0, $zero, 161   d
		 7'b0011110: Instruct<=32'b101011_00000_01000_0000000000110100; //sw    $t0, 52($zero)
		 7'b0011111: Instruct<=32'b001001_00000_01000_0000000010000110; //addiu $t0, $zero, 134   e
		 7'b0100000: Instruct<=32'b101011_00000_01000_0000000000111000; //sw    $t0, 56($zero)
		 7'b0100001: Instruct<=32'b001001_00000_01000_0000000010001110; //addiu $t0, $zero, 142   f
		 7'b0100010: Instruct<=32'b101011_00000_01000_0000000000111100; //sw    $t0, 60($zero)
		 //Initial v0=1
		 7'b0100011: Instruct<=32'b001001_00000_00010_0000000000000001; //addiu $v0, $zero, 1       //$v0:AN
		 //record the two 8bits numbers
		 7'b0100100: Instruct<=32'b000000_00000_00000_0000000000000000;   //nop
		 7'b0100101: Instruct<=32'b100011_10000_10001_0000000000011100;   //lw   $s1, 28($s0)        //$s1:UART_RXD
		 7'b0100110: Instruct<=32'b000000_00000_10001_01001_00000_100000; //add  $t1, $s1, $zero
		 7'b0100111: Instruct<=32'b100011_10000_10010_0000000000011100;   //lw   $s2, 28($s0)        //$s2:UART_RXD
		 7'b0101000: Instruct<=32'b000000_00000_10010_01010_00000_100000; //add  $t2, $s2, $zero
		 7'b0101001: Instruct<=32'b000100_01001_00000_0000000000001000;   //beq  $t1, $zero, caseC   //num1==0,result=num2
		 7'b0101010: Instruct<=32'b000100_01010_00000_0000000000001001;   //beq  $t2, $zero, caseD   //num2==0,result=num1
	  	//Loop1:
		 7'b0101011: Instruct<=32'b000100_01001_01010_0000000000001000;   //beq  $t1, $t2, caseD
		 7'b0101100: Instruct<=32'b000000_01001_01010_01000_00000_101010; //slt  $t0, $t1, $t2
		 7'b0101101: Instruct<=32'b000101_01000_00000_0000000000000010;   //bne  $t0, $zero, caseB
		 //caseA:
		 7'b0101110: Instruct<=32'b000000_01001_01010_01001_00000_100010; //sub  $t1, $t1, $t2       //num1>num2
		 7'b0101111: Instruct<=32'b000010_00000000000000000000101011;     //j    Loop1
		 //caseB:
		 7'b0110000: Instruct<=32'b000000_01010_01001_01010_00000_100010; //sub  $t2, $t2, $t1       //num2>num1
		 7'b0110001: Instruct<=32'b000010_00000000000000000000101011;     //j    Loop1
		 //caseC:
		 7'b0110010: Instruct<=32'b000000_01010_00000_00011_00000_100000; //add  $v1, $t2, $zero     //$v1:result
		 7'b0110011: Instruct<=32'b000010_00000000000000000000110101;     //j    AN                  
	  	//caseD:                  
		 7'b0110100: Instruct<=32'b000000_01010_00000_00011_00000_100000; //add  $v1, $t2, $zero     	 
		 //AN:           
		 7'b0110101: Instruct<=32'b000000_00000_00010_01011_00001_000010; //srl  $t3, $v0, 1         
		 7'b0110110: Instruct<=32'b000100_01011_00000_0000000000001000;   //beq  $t3, $zero, num1     //digital:num1
		 7'b0110111: Instruct<=32'b000000_00000_00010_01011_00010_000010; //srl  $t3, $v0, 2
		 7'b0111000: Instruct<=32'b000100_01011_00000_0000000000001001;   //beq  $t3, $zero, num2     //digital:num2
		 7'b0111001: Instruct<=32'b000000_00000_00010_01011_00011_000010; //srl  $t3, $v0, 3         
		 7'b0111010: Instruct<=32'b000100_01011_00000_0000000000001010;   //beq  $t3, $zero, num3     //digital:num3
     7'b0111011: Instruct<=32'b001001_00000_00010_0000000000000001;   //addiu $v0, $zero, 1       //digital:num4
 		 7'b0111100: Instruct<=32'b000000_00000_10010_10011_00100_000010; //srl  $s3, $s2, 4		 
		 7'b0111101: Instruct<=32'b000000_00000_10011_10011_00010_000000; //sll  $s3, $s3, 2
		 7'b0111110: Instruct<=32'b000010_00000000000000000001001001;     //j     Output
		 //num1:
		 7'b0111111: Instruct<=32'b001100_10001_10011_0000000000001111;   //andi $s3, $s1, 15 
		 7'b1000000: Instruct<=32'b000000_00000_10011_10011_00010_000000; //sll  $s3, $s3, 2 
		 7'b1000001: Instruct<=32'b000010_00000000000000000001001000;     //j    shift 
		 //num2:
		 7'b1000010: Instruct<=32'b000000_00000_10001_10011_00100_000010; //srl  $s3, $s1, 4		 
		 7'b1000011: Instruct<=32'b000000_00000_10011_10011_00010_000000; //sll  $s3, $s3, 2
		 7'b1000100: Instruct<=32'b000010_00000000000000000001001000;     //j    shift
		 //num3:
		 7'b1000101: Instruct<=32'b001100_10010_10011_0000000000001111;   //andi $s3, $s2, 15 
		 7'b1000110: Instruct<=32'b000000_00000_10011_10011_00010_000000; //sll  $s3, $s3, 2 
		 7'b1000111: Instruct<=32'b000010_00000000000000000001001000;     //j    shift 		 
		 //shift:
		 7'b1001000: Instruct<=32'b000000_00000_00010_00010_00001_000000; //sll  $v0, $v0, 1
		 //Output:
		 7'b1001001: Instruct<=32'b000010_00000000000000000001001001;     //j   Output
		 7'b1001010: Instruct<=32'b00000000000000000000000000000000;      //nop
		 7'b1001011: Instruct<=32'b00000000000000000000000000000000;      //nop
		 7'b1001100: Instruct<=32'b000010_00000000000000000000100100;     //j   preparation
	  	//reset:
		 7'b1001101: Instruct<=32'b001001_00000_10100_0000000000000011;   //addiu $s4, $zero, 3  //$s4:TCON=3
		 7'b1001110: Instruct<=32'b001111_00000_10000_0100000000000000;   //lui   $s0, 16384
		 7'b1001111: Instruct<=32'b101011_10000_10100_0000000000001000;   //sw    $s4, 8($s0)
     7'b1010000: Instruct<=32'b001001_00000_10111_0000000000000011;   //addiu $s7, $zero, 3  
     7'b1010001: Instruct<=32'b000000_00000_10111_10111_00010_000000; //sll   $s7, $s7, 2 
		 7'b1010010: Instruct<=32'b000000_10111_00000_00000_00000_001000; //jr    $s7
		 //ILLOP:
		 7'b1010011: Instruct<=32'b101011_10000_10100_0000000000001000;   //sw   $s4, 8($s0)
		 7'b1010100: Instruct<=32'b100011_10011_10101_0000000000000000;   //lw   $s5, 0($s3)     
		 7'b1010101: Instruct<=32'b000000_00000_00010_10110_01000_000000; //sll  $s6, $v0, 8     //$s6:{AN,digital}
		 7'b1010110: Instruct<=32'b000000_10101_10110_10110_00000_100000; //add  $s6, $s5, $s6
	   7'b1010111: Instruct<=32'b101011_10000_10110_0000000000010100;   //sw   $s6, 20($s0)
     7'b1011000: Instruct<=32'b101011_10000_00011_0000000000001100;   //sw   $v1, 12($s0)
     7'b1011001: Instruct<=32'b101011_10000_00011_0000000000011000;   //sw   $v1, 24($s0)
		 7'b1011010: Instruct<=32'b000000_11010_00000_00000_00000_001000; //jr   $xp
		 default:	Instruct<=32'b0;
		endcase
	 end
 end

endmodule
